VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_sram_1r1w_128x512_128
   CLASS BLOCK ;
   SIZE 1250.9 BY 641.62 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  161.16 0.0 161.54 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  167.28 0.0 167.66 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  173.4 0.0 173.78 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  178.84 0.0 179.22 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  184.96 0.0 185.34 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  191.08 0.0 191.46 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  196.52 0.0 196.9 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  202.64 0.0 203.02 1.06 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  208.08 0.0 208.46 1.06 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  214.2 0.0 214.58 1.06 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  220.32 0.0 220.7 1.06 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  225.76 0.0 226.14 1.06 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  231.88 0.0 232.26 1.06 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  237.32 0.0 237.7 1.06 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  243.44 0.0 243.82 1.06 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  249.56 0.0 249.94 1.06 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  255.0 0.0 255.38 1.06 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  261.12 0.0 261.5 1.06 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  266.56 0.0 266.94 1.06 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  272.68 0.0 273.06 1.06 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  278.12 0.0 278.5 1.06 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  284.24 0.0 284.62 1.06 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  289.68 0.0 290.06 1.06 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  295.8 0.0 296.18 1.06 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  301.92 0.0 302.3 1.06 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  307.36 0.0 307.74 1.06 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  313.48 0.0 313.86 1.06 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  319.6 0.0 319.98 1.06 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  325.04 0.0 325.42 1.06 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  331.16 0.0 331.54 1.06 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  336.6 0.0 336.98 1.06 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  342.72 0.0 343.1 1.06 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  348.84 0.0 349.22 1.06 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  354.28 0.0 354.66 1.06 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  360.4 0.0 360.78 1.06 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  365.84 0.0 366.22 1.06 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  371.96 0.0 372.34 1.06 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  378.08 0.0 378.46 1.06 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  383.52 0.0 383.9 1.06 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  388.96 0.0 389.34 1.06 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  395.08 0.0 395.46 1.06 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  400.52 0.0 400.9 1.06 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  406.64 0.0 407.02 1.06 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  412.76 0.0 413.14 1.06 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  418.2 0.0 418.58 1.06 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  424.32 0.0 424.7 1.06 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  429.76 0.0 430.14 1.06 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  435.88 0.0 436.26 1.06 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  442.0 0.0 442.38 1.06 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  447.44 0.0 447.82 1.06 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  453.56 0.0 453.94 1.06 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  459.68 0.0 460.06 1.06 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  465.12 0.0 465.5 1.06 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  471.24 0.0 471.62 1.06 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  476.68 0.0 477.06 1.06 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  482.8 0.0 483.18 1.06 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  488.24 0.0 488.62 1.06 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  494.36 0.0 494.74 1.06 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  500.48 0.0 500.86 1.06 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  505.92 0.0 506.3 1.06 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  512.04 0.0 512.42 1.06 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  518.16 0.0 518.54 1.06 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  523.6 0.0 523.98 1.06 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  529.72 0.0 530.1 1.06 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  535.16 0.0 535.54 1.06 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  541.28 0.0 541.66 1.06 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  546.72 0.0 547.1 1.06 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  552.84 0.0 553.22 1.06 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  558.28 0.0 558.66 1.06 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  564.4 0.0 564.78 1.06 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  570.52 0.0 570.9 1.06 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  576.64 0.0 577.02 1.06 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  582.08 0.0 582.46 1.06 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  587.52 0.0 587.9 1.06 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  593.64 0.0 594.02 1.06 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  599.76 0.0 600.14 1.06 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  605.2 0.0 605.58 1.06 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  611.32 0.0 611.7 1.06 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  616.76 0.0 617.14 1.06 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  622.88 0.0 623.26 1.06 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  628.32 0.0 628.7 1.06 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  634.44 0.0 634.82 1.06 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  640.56 0.0 640.94 1.06 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  646.68 0.0 647.06 1.06 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  652.12 0.0 652.5 1.06 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  658.24 0.0 658.62 1.06 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  663.68 0.0 664.06 1.06 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  669.8 0.0 670.18 1.06 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  675.24 0.0 675.62 1.06 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  681.36 0.0 681.74 1.06 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  686.8 0.0 687.18 1.06 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  692.92 0.0 693.3 1.06 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  698.36 0.0 698.74 1.06 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  704.48 0.0 704.86 1.06 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  710.6 0.0 710.98 1.06 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  716.04 0.0 716.42 1.06 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  722.16 0.0 722.54 1.06 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  727.6 0.0 727.98 1.06 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  733.72 0.0 734.1 1.06 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  739.84 0.0 740.22 1.06 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  745.96 0.0 746.34 1.06 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  751.4 0.0 751.78 1.06 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  757.52 0.0 757.9 1.06 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  762.96 0.0 763.34 1.06 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  769.08 0.0 769.46 1.06 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  775.2 0.0 775.58 1.06 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  780.64 0.0 781.02 1.06 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  786.08 0.0 786.46 1.06 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  792.2 0.0 792.58 1.06 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  798.32 0.0 798.7 1.06 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  803.76 0.0 804.14 1.06 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  809.88 0.0 810.26 1.06 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  816.0 0.0 816.38 1.06 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  821.44 0.0 821.82 1.06 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  827.56 0.0 827.94 1.06 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  833.0 0.0 833.38 1.06 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  839.12 0.0 839.5 1.06 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  845.24 0.0 845.62 1.06 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  850.68 0.0 851.06 1.06 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  856.12 0.0 856.5 1.06 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  862.24 0.0 862.62 1.06 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  868.36 0.0 868.74 1.06 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  874.48 0.0 874.86 1.06 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  879.92 0.0 880.3 1.06 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  886.04 0.0 886.42 1.06 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  891.48 0.0 891.86 1.06 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  896.92 0.0 897.3 1.06 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  903.04 0.0 903.42 1.06 ;
      END
   END din0[127]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  155.72 0.0 156.1 1.06 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  144.16 0.0 144.54 1.06 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  144.84 0.0 145.22 1.06 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  142.12 0.0 142.5 1.06 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 148.92 1.06 149.3 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 154.36 1.06 154.74 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 163.2 1.06 163.58 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 167.96 1.06 168.34 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 176.8 1.06 177.18 ;
      END
   END addr0[8]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1088.0 640.56 1088.38 641.62 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1109.08 0.0 1109.46 1.06 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1102.96 0.0 1103.34 1.06 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1103.64 0.0 1104.02 1.06 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1108.4 0.0 1108.78 1.06 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1107.72 0.0 1108.1 1.06 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1104.32 0.0 1104.7 1.06 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1105.0 0.0 1105.38 1.06 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1105.68 0.0 1106.06 1.06 ;
      END
   END addr1[8]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 24.48 1.06 24.86 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1249.84 625.6 1250.9 625.98 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  30.6 0.0 30.98 1.06 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1219.24 640.56 1219.62 641.62 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  225.76 640.56 226.14 641.62 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  232.56 640.56 232.94 641.62 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  238.68 640.56 239.06 641.62 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  244.12 640.56 244.5 641.62 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  250.92 640.56 251.3 641.62 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  257.04 640.56 257.42 641.62 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  263.16 640.56 263.54 641.62 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  269.96 640.56 270.34 641.62 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  275.4 640.56 275.78 641.62 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  282.88 640.56 283.26 641.62 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  289.0 640.56 289.38 641.62 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  295.12 640.56 295.5 641.62 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  300.56 640.56 300.94 641.62 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  307.36 640.56 307.74 641.62 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  313.48 640.56 313.86 641.62 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  319.6 640.56 319.98 641.62 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  325.72 640.56 326.1 641.62 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  332.52 640.56 332.9 641.62 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  337.96 640.56 338.34 641.62 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  344.08 640.56 344.46 641.62 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  350.88 640.56 351.26 641.62 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  357.68 640.56 358.06 641.62 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  363.12 640.56 363.5 641.62 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  369.24 640.56 369.62 641.62 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  376.04 640.56 376.42 641.62 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  382.16 640.56 382.54 641.62 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  387.6 640.56 387.98 641.62 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  394.4 640.56 394.78 641.62 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  400.52 640.56 400.9 641.62 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  407.32 640.56 407.7 641.62 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  413.44 640.56 413.82 641.62 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  418.88 640.56 419.26 641.62 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  426.36 640.56 426.74 641.62 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  432.48 640.56 432.86 641.62 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  438.6 640.56 438.98 641.62 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  444.04 640.56 444.42 641.62 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  450.16 640.56 450.54 641.62 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  456.28 640.56 456.66 641.62 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  463.08 640.56 463.46 641.62 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  469.88 640.56 470.26 641.62 ;
      END
   END dout1[39]
   PIN dout1[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  475.32 640.56 475.7 641.62 ;
      END
   END dout1[40]
   PIN dout1[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  481.44 640.56 481.82 641.62 ;
      END
   END dout1[41]
   PIN dout1[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  487.56 640.56 487.94 641.62 ;
      END
   END dout1[42]
   PIN dout1[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  494.36 640.56 494.74 641.62 ;
      END
   END dout1[43]
   PIN dout1[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  500.48 640.56 500.86 641.62 ;
      END
   END dout1[44]
   PIN dout1[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  507.28 640.56 507.66 641.62 ;
      END
   END dout1[45]
   PIN dout1[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  513.4 640.56 513.78 641.62 ;
      END
   END dout1[46]
   PIN dout1[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  518.84 640.56 519.22 641.62 ;
      END
   END dout1[47]
   PIN dout1[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  525.64 640.56 526.02 641.62 ;
      END
   END dout1[48]
   PIN dout1[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  531.76 640.56 532.14 641.62 ;
      END
   END dout1[49]
   PIN dout1[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  538.56 640.56 538.94 641.62 ;
      END
   END dout1[50]
   PIN dout1[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  544.0 640.56 544.38 641.62 ;
      END
   END dout1[51]
   PIN dout1[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  550.8 640.56 551.18 641.62 ;
      END
   END dout1[52]
   PIN dout1[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  556.24 640.56 556.62 641.62 ;
      END
   END dout1[53]
   PIN dout1[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  563.04 640.56 563.42 641.62 ;
      END
   END dout1[54]
   PIN dout1[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  568.48 640.56 568.86 641.62 ;
      END
   END dout1[55]
   PIN dout1[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  575.28 640.56 575.66 641.62 ;
      END
   END dout1[56]
   PIN dout1[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  582.08 640.56 582.46 641.62 ;
      END
   END dout1[57]
   PIN dout1[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  587.52 640.56 587.9 641.62 ;
      END
   END dout1[58]
   PIN dout1[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  593.64 640.56 594.02 641.62 ;
      END
   END dout1[59]
   PIN dout1[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  601.12 640.56 601.5 641.62 ;
      END
   END dout1[60]
   PIN dout1[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  607.24 640.56 607.62 641.62 ;
      END
   END dout1[61]
   PIN dout1[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  612.68 640.56 613.06 641.62 ;
      END
   END dout1[62]
   PIN dout1[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  618.8 640.56 619.18 641.62 ;
      END
   END dout1[63]
   PIN dout1[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  624.92 640.56 625.3 641.62 ;
      END
   END dout1[64]
   PIN dout1[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  631.04 640.56 631.42 641.62 ;
      END
   END dout1[65]
   PIN dout1[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  637.16 640.56 637.54 641.62 ;
      END
   END dout1[66]
   PIN dout1[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  643.96 640.56 644.34 641.62 ;
      END
   END dout1[67]
   PIN dout1[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  650.76 640.56 651.14 641.62 ;
      END
   END dout1[68]
   PIN dout1[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  656.88 640.56 657.26 641.62 ;
      END
   END dout1[69]
   PIN dout1[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  662.32 640.56 662.7 641.62 ;
      END
   END dout1[70]
   PIN dout1[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  669.12 640.56 669.5 641.62 ;
      END
   END dout1[71]
   PIN dout1[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  675.92 640.56 676.3 641.62 ;
      END
   END dout1[72]
   PIN dout1[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  682.04 640.56 682.42 641.62 ;
      END
   END dout1[73]
   PIN dout1[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  687.48 640.56 687.86 641.62 ;
      END
   END dout1[74]
   PIN dout1[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  693.6 640.56 693.98 641.62 ;
      END
   END dout1[75]
   PIN dout1[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  700.4 640.56 700.78 641.62 ;
      END
   END dout1[76]
   PIN dout1[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  707.2 640.56 707.58 641.62 ;
      END
   END dout1[77]
   PIN dout1[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  712.64 640.56 713.02 641.62 ;
      END
   END dout1[78]
   PIN dout1[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  719.44 640.56 719.82 641.62 ;
      END
   END dout1[79]
   PIN dout1[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  725.56 640.56 725.94 641.62 ;
      END
   END dout1[80]
   PIN dout1[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  731.0 640.56 731.38 641.62 ;
      END
   END dout1[81]
   PIN dout1[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  737.12 640.56 737.5 641.62 ;
      END
   END dout1[82]
   PIN dout1[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  743.92 640.56 744.3 641.62 ;
      END
   END dout1[83]
   PIN dout1[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  750.72 640.56 751.1 641.62 ;
      END
   END dout1[84]
   PIN dout1[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  756.16 640.56 756.54 641.62 ;
      END
   END dout1[85]
   PIN dout1[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  762.28 640.56 762.66 641.62 ;
      END
   END dout1[86]
   PIN dout1[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  769.08 640.56 769.46 641.62 ;
      END
   END dout1[87]
   PIN dout1[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  775.2 640.56 775.58 641.62 ;
      END
   END dout1[88]
   PIN dout1[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  780.64 640.56 781.02 641.62 ;
      END
   END dout1[89]
   PIN dout1[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  787.44 640.56 787.82 641.62 ;
      END
   END dout1[90]
   PIN dout1[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  793.56 640.56 793.94 641.62 ;
      END
   END dout1[91]
   PIN dout1[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  800.36 640.56 800.74 641.62 ;
      END
   END dout1[92]
   PIN dout1[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  805.8 640.56 806.18 641.62 ;
      END
   END dout1[93]
   PIN dout1[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  812.6 640.56 812.98 641.62 ;
      END
   END dout1[94]
   PIN dout1[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  819.4 640.56 819.78 641.62 ;
      END
   END dout1[95]
   PIN dout1[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  825.52 640.56 825.9 641.62 ;
      END
   END dout1[96]
   PIN dout1[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  830.96 640.56 831.34 641.62 ;
      END
   END dout1[97]
   PIN dout1[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  837.76 640.56 838.14 641.62 ;
      END
   END dout1[98]
   PIN dout1[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  843.2 640.56 843.58 641.62 ;
      END
   END dout1[99]
   PIN dout1[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  849.32 640.56 849.7 641.62 ;
      END
   END dout1[100]
   PIN dout1[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  856.12 640.56 856.5 641.62 ;
      END
   END dout1[101]
   PIN dout1[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  862.92 640.56 863.3 641.62 ;
      END
   END dout1[102]
   PIN dout1[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  868.36 640.56 868.74 641.62 ;
      END
   END dout1[103]
   PIN dout1[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  874.48 640.56 874.86 641.62 ;
      END
   END dout1[104]
   PIN dout1[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  880.6 640.56 880.98 641.62 ;
      END
   END dout1[105]
   PIN dout1[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  887.4 640.56 887.78 641.62 ;
      END
   END dout1[106]
   PIN dout1[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  894.2 640.56 894.58 641.62 ;
      END
   END dout1[107]
   PIN dout1[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  900.32 640.56 900.7 641.62 ;
      END
   END dout1[108]
   PIN dout1[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  905.76 640.56 906.14 641.62 ;
      END
   END dout1[109]
   PIN dout1[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  911.88 640.56 912.26 641.62 ;
      END
   END dout1[110]
   PIN dout1[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  918.68 640.56 919.06 641.62 ;
      END
   END dout1[111]
   PIN dout1[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  924.8 640.56 925.18 641.62 ;
      END
   END dout1[112]
   PIN dout1[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  931.6 640.56 931.98 641.62 ;
      END
   END dout1[113]
   PIN dout1[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  937.04 640.56 937.42 641.62 ;
      END
   END dout1[114]
   PIN dout1[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  943.16 640.56 943.54 641.62 ;
      END
   END dout1[115]
   PIN dout1[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  949.96 640.56 950.34 641.62 ;
      END
   END dout1[116]
   PIN dout1[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  955.4 640.56 955.78 641.62 ;
      END
   END dout1[117]
   PIN dout1[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  962.2 640.56 962.58 641.62 ;
      END
   END dout1[118]
   PIN dout1[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  969.0 640.56 969.38 641.62 ;
      END
   END dout1[119]
   PIN dout1[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  974.44 640.56 974.82 641.62 ;
      END
   END dout1[120]
   PIN dout1[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  980.56 640.56 980.94 641.62 ;
      END
   END dout1[121]
   PIN dout1[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  987.36 640.56 987.74 641.62 ;
      END
   END dout1[122]
   PIN dout1[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  994.16 640.56 994.54 641.62 ;
      END
   END dout1[123]
   PIN dout1[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  999.6 640.56 999.98 641.62 ;
      END
   END dout1[124]
   PIN dout1[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1005.72 640.56 1006.1 641.62 ;
      END
   END dout1[125]
   PIN dout1[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1012.52 640.56 1012.9 641.62 ;
      END
   END dout1[126]
   PIN dout1[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1018.64 640.56 1019.02 641.62 ;
      END
   END dout1[127]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  1245.76 3.4 1247.5 638.22 ;
         LAYER met3 ;
         RECT  3.4 3.4 1247.5 5.14 ;
         LAYER met4 ;
         RECT  3.4 3.4 5.14 638.22 ;
         LAYER met3 ;
         RECT  3.4 636.48 1247.5 638.22 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  0.0 0.0 1250.9 1.74 ;
         LAYER met3 ;
         RECT  0.0 639.88 1250.9 641.62 ;
         LAYER met4 ;
         RECT  1249.16 0.0 1250.9 641.62 ;
         LAYER met4 ;
         RECT  0.0 0.0 1.74 641.62 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 1250.28 641.0 ;
   LAYER  met2 ;
      RECT  0.62 0.62 1250.28 641.0 ;
   LAYER  met3 ;
      RECT  1.66 148.32 1250.28 149.9 ;
      RECT  0.62 149.9 1.66 153.76 ;
      RECT  0.62 155.34 1.66 162.6 ;
      RECT  0.62 164.18 1.66 167.36 ;
      RECT  0.62 168.94 1.66 176.2 ;
      RECT  0.62 25.46 1.66 148.32 ;
      RECT  1.66 149.9 1249.24 625.0 ;
      RECT  1.66 625.0 1249.24 626.58 ;
      RECT  1249.24 149.9 1250.28 625.0 ;
      RECT  1.66 2.8 2.8 5.74 ;
      RECT  1.66 5.74 2.8 148.32 ;
      RECT  2.8 5.74 1248.1 148.32 ;
      RECT  1248.1 2.8 1250.28 5.74 ;
      RECT  1248.1 5.74 1250.28 148.32 ;
      RECT  1.66 626.58 2.8 635.88 ;
      RECT  1.66 635.88 2.8 638.82 ;
      RECT  2.8 626.58 1248.1 635.88 ;
      RECT  1248.1 626.58 1249.24 635.88 ;
      RECT  1248.1 635.88 1249.24 638.82 ;
      RECT  0.62 2.34 1.66 23.88 ;
      RECT  1.66 2.34 2.8 2.8 ;
      RECT  2.8 2.34 1248.1 2.8 ;
      RECT  1248.1 2.34 1250.28 2.8 ;
      RECT  0.62 177.78 1.66 639.28 ;
      RECT  1249.24 626.58 1250.28 639.28 ;
      RECT  1.66 638.82 2.8 639.28 ;
      RECT  2.8 638.82 1248.1 639.28 ;
      RECT  1248.1 638.82 1249.24 639.28 ;
   LAYER  met4 ;
      RECT  160.56 1.66 162.14 641.0 ;
      RECT  162.14 0.62 166.68 1.66 ;
      RECT  168.26 0.62 172.8 1.66 ;
      RECT  174.38 0.62 178.24 1.66 ;
      RECT  179.82 0.62 184.36 1.66 ;
      RECT  185.94 0.62 190.48 1.66 ;
      RECT  192.06 0.62 195.92 1.66 ;
      RECT  197.5 0.62 202.04 1.66 ;
      RECT  203.62 0.62 207.48 1.66 ;
      RECT  209.06 0.62 213.6 1.66 ;
      RECT  215.18 0.62 219.72 1.66 ;
      RECT  221.3 0.62 225.16 1.66 ;
      RECT  226.74 0.62 231.28 1.66 ;
      RECT  232.86 0.62 236.72 1.66 ;
      RECT  238.3 0.62 242.84 1.66 ;
      RECT  244.42 0.62 248.96 1.66 ;
      RECT  250.54 0.62 254.4 1.66 ;
      RECT  255.98 0.62 260.52 1.66 ;
      RECT  262.1 0.62 265.96 1.66 ;
      RECT  267.54 0.62 272.08 1.66 ;
      RECT  273.66 0.62 277.52 1.66 ;
      RECT  279.1 0.62 283.64 1.66 ;
      RECT  285.22 0.62 289.08 1.66 ;
      RECT  290.66 0.62 295.2 1.66 ;
      RECT  296.78 0.62 301.32 1.66 ;
      RECT  302.9 0.62 306.76 1.66 ;
      RECT  308.34 0.62 312.88 1.66 ;
      RECT  314.46 0.62 319.0 1.66 ;
      RECT  320.58 0.62 324.44 1.66 ;
      RECT  326.02 0.62 330.56 1.66 ;
      RECT  332.14 0.62 336.0 1.66 ;
      RECT  337.58 0.62 342.12 1.66 ;
      RECT  343.7 0.62 348.24 1.66 ;
      RECT  349.82 0.62 353.68 1.66 ;
      RECT  355.26 0.62 359.8 1.66 ;
      RECT  361.38 0.62 365.24 1.66 ;
      RECT  366.82 0.62 371.36 1.66 ;
      RECT  372.94 0.62 377.48 1.66 ;
      RECT  379.06 0.62 382.92 1.66 ;
      RECT  384.5 0.62 388.36 1.66 ;
      RECT  389.94 0.62 394.48 1.66 ;
      RECT  396.06 0.62 399.92 1.66 ;
      RECT  401.5 0.62 406.04 1.66 ;
      RECT  407.62 0.62 412.16 1.66 ;
      RECT  413.74 0.62 417.6 1.66 ;
      RECT  419.18 0.62 423.72 1.66 ;
      RECT  425.3 0.62 429.16 1.66 ;
      RECT  430.74 0.62 435.28 1.66 ;
      RECT  436.86 0.62 441.4 1.66 ;
      RECT  442.98 0.62 446.84 1.66 ;
      RECT  448.42 0.62 452.96 1.66 ;
      RECT  454.54 0.62 459.08 1.66 ;
      RECT  460.66 0.62 464.52 1.66 ;
      RECT  466.1 0.62 470.64 1.66 ;
      RECT  472.22 0.62 476.08 1.66 ;
      RECT  477.66 0.62 482.2 1.66 ;
      RECT  483.78 0.62 487.64 1.66 ;
      RECT  489.22 0.62 493.76 1.66 ;
      RECT  495.34 0.62 499.88 1.66 ;
      RECT  501.46 0.62 505.32 1.66 ;
      RECT  506.9 0.62 511.44 1.66 ;
      RECT  513.02 0.62 517.56 1.66 ;
      RECT  519.14 0.62 523.0 1.66 ;
      RECT  524.58 0.62 529.12 1.66 ;
      RECT  530.7 0.62 534.56 1.66 ;
      RECT  536.14 0.62 540.68 1.66 ;
      RECT  542.26 0.62 546.12 1.66 ;
      RECT  547.7 0.62 552.24 1.66 ;
      RECT  553.82 0.62 557.68 1.66 ;
      RECT  559.26 0.62 563.8 1.66 ;
      RECT  565.38 0.62 569.92 1.66 ;
      RECT  571.5 0.62 576.04 1.66 ;
      RECT  577.62 0.62 581.48 1.66 ;
      RECT  583.06 0.62 586.92 1.66 ;
      RECT  588.5 0.62 593.04 1.66 ;
      RECT  594.62 0.62 599.16 1.66 ;
      RECT  600.74 0.62 604.6 1.66 ;
      RECT  606.18 0.62 610.72 1.66 ;
      RECT  612.3 0.62 616.16 1.66 ;
      RECT  617.74 0.62 622.28 1.66 ;
      RECT  623.86 0.62 627.72 1.66 ;
      RECT  629.3 0.62 633.84 1.66 ;
      RECT  635.42 0.62 639.96 1.66 ;
      RECT  641.54 0.62 646.08 1.66 ;
      RECT  647.66 0.62 651.52 1.66 ;
      RECT  653.1 0.62 657.64 1.66 ;
      RECT  659.22 0.62 663.08 1.66 ;
      RECT  664.66 0.62 669.2 1.66 ;
      RECT  670.78 0.62 674.64 1.66 ;
      RECT  676.22 0.62 680.76 1.66 ;
      RECT  682.34 0.62 686.2 1.66 ;
      RECT  687.78 0.62 692.32 1.66 ;
      RECT  693.9 0.62 697.76 1.66 ;
      RECT  699.34 0.62 703.88 1.66 ;
      RECT  705.46 0.62 710.0 1.66 ;
      RECT  711.58 0.62 715.44 1.66 ;
      RECT  717.02 0.62 721.56 1.66 ;
      RECT  723.14 0.62 727.0 1.66 ;
      RECT  728.58 0.62 733.12 1.66 ;
      RECT  734.7 0.62 739.24 1.66 ;
      RECT  740.82 0.62 745.36 1.66 ;
      RECT  746.94 0.62 750.8 1.66 ;
      RECT  752.38 0.62 756.92 1.66 ;
      RECT  758.5 0.62 762.36 1.66 ;
      RECT  763.94 0.62 768.48 1.66 ;
      RECT  770.06 0.62 774.6 1.66 ;
      RECT  776.18 0.62 780.04 1.66 ;
      RECT  781.62 0.62 785.48 1.66 ;
      RECT  787.06 0.62 791.6 1.66 ;
      RECT  793.18 0.62 797.72 1.66 ;
      RECT  799.3 0.62 803.16 1.66 ;
      RECT  804.74 0.62 809.28 1.66 ;
      RECT  810.86 0.62 815.4 1.66 ;
      RECT  816.98 0.62 820.84 1.66 ;
      RECT  822.42 0.62 826.96 1.66 ;
      RECT  828.54 0.62 832.4 1.66 ;
      RECT  833.98 0.62 838.52 1.66 ;
      RECT  840.1 0.62 844.64 1.66 ;
      RECT  846.22 0.62 850.08 1.66 ;
      RECT  851.66 0.62 855.52 1.66 ;
      RECT  857.1 0.62 861.64 1.66 ;
      RECT  863.22 0.62 867.76 1.66 ;
      RECT  869.34 0.62 873.88 1.66 ;
      RECT  875.46 0.62 879.32 1.66 ;
      RECT  880.9 0.62 885.44 1.66 ;
      RECT  887.02 0.62 890.88 1.66 ;
      RECT  892.46 0.62 896.32 1.66 ;
      RECT  897.9 0.62 902.44 1.66 ;
      RECT  156.7 0.62 160.56 1.66 ;
      RECT  145.82 0.62 155.12 1.66 ;
      RECT  143.1 0.62 143.56 1.66 ;
      RECT  162.14 1.66 1087.4 639.96 ;
      RECT  1087.4 1.66 1088.98 639.96 ;
      RECT  904.02 0.62 1102.36 1.66 ;
      RECT  1106.66 0.62 1107.12 1.66 ;
      RECT  31.58 0.62 141.52 1.66 ;
      RECT  1088.98 639.96 1218.64 641.0 ;
      RECT  162.14 639.96 225.16 641.0 ;
      RECT  226.74 639.96 231.96 641.0 ;
      RECT  233.54 639.96 238.08 641.0 ;
      RECT  239.66 639.96 243.52 641.0 ;
      RECT  245.1 639.96 250.32 641.0 ;
      RECT  251.9 639.96 256.44 641.0 ;
      RECT  258.02 639.96 262.56 641.0 ;
      RECT  264.14 639.96 269.36 641.0 ;
      RECT  270.94 639.96 274.8 641.0 ;
      RECT  276.38 639.96 282.28 641.0 ;
      RECT  283.86 639.96 288.4 641.0 ;
      RECT  289.98 639.96 294.52 641.0 ;
      RECT  296.1 639.96 299.96 641.0 ;
      RECT  301.54 639.96 306.76 641.0 ;
      RECT  308.34 639.96 312.88 641.0 ;
      RECT  314.46 639.96 319.0 641.0 ;
      RECT  320.58 639.96 325.12 641.0 ;
      RECT  326.7 639.96 331.92 641.0 ;
      RECT  333.5 639.96 337.36 641.0 ;
      RECT  338.94 639.96 343.48 641.0 ;
      RECT  345.06 639.96 350.28 641.0 ;
      RECT  351.86 639.96 357.08 641.0 ;
      RECT  358.66 639.96 362.52 641.0 ;
      RECT  364.1 639.96 368.64 641.0 ;
      RECT  370.22 639.96 375.44 641.0 ;
      RECT  377.02 639.96 381.56 641.0 ;
      RECT  383.14 639.96 387.0 641.0 ;
      RECT  388.58 639.96 393.8 641.0 ;
      RECT  395.38 639.96 399.92 641.0 ;
      RECT  401.5 639.96 406.72 641.0 ;
      RECT  408.3 639.96 412.84 641.0 ;
      RECT  414.42 639.96 418.28 641.0 ;
      RECT  419.86 639.96 425.76 641.0 ;
      RECT  427.34 639.96 431.88 641.0 ;
      RECT  433.46 639.96 438.0 641.0 ;
      RECT  439.58 639.96 443.44 641.0 ;
      RECT  445.02 639.96 449.56 641.0 ;
      RECT  451.14 639.96 455.68 641.0 ;
      RECT  457.26 639.96 462.48 641.0 ;
      RECT  464.06 639.96 469.28 641.0 ;
      RECT  470.86 639.96 474.72 641.0 ;
      RECT  476.3 639.96 480.84 641.0 ;
      RECT  482.42 639.96 486.96 641.0 ;
      RECT  488.54 639.96 493.76 641.0 ;
      RECT  495.34 639.96 499.88 641.0 ;
      RECT  501.46 639.96 506.68 641.0 ;
      RECT  508.26 639.96 512.8 641.0 ;
      RECT  514.38 639.96 518.24 641.0 ;
      RECT  519.82 639.96 525.04 641.0 ;
      RECT  526.62 639.96 531.16 641.0 ;
      RECT  532.74 639.96 537.96 641.0 ;
      RECT  539.54 639.96 543.4 641.0 ;
      RECT  544.98 639.96 550.2 641.0 ;
      RECT  551.78 639.96 555.64 641.0 ;
      RECT  557.22 639.96 562.44 641.0 ;
      RECT  564.02 639.96 567.88 641.0 ;
      RECT  569.46 639.96 574.68 641.0 ;
      RECT  576.26 639.96 581.48 641.0 ;
      RECT  583.06 639.96 586.92 641.0 ;
      RECT  588.5 639.96 593.04 641.0 ;
      RECT  594.62 639.96 600.52 641.0 ;
      RECT  602.1 639.96 606.64 641.0 ;
      RECT  608.22 639.96 612.08 641.0 ;
      RECT  613.66 639.96 618.2 641.0 ;
      RECT  619.78 639.96 624.32 641.0 ;
      RECT  625.9 639.96 630.44 641.0 ;
      RECT  632.02 639.96 636.56 641.0 ;
      RECT  638.14 639.96 643.36 641.0 ;
      RECT  644.94 639.96 650.16 641.0 ;
      RECT  651.74 639.96 656.28 641.0 ;
      RECT  657.86 639.96 661.72 641.0 ;
      RECT  663.3 639.96 668.52 641.0 ;
      RECT  670.1 639.96 675.32 641.0 ;
      RECT  676.9 639.96 681.44 641.0 ;
      RECT  683.02 639.96 686.88 641.0 ;
      RECT  688.46 639.96 693.0 641.0 ;
      RECT  694.58 639.96 699.8 641.0 ;
      RECT  701.38 639.96 706.6 641.0 ;
      RECT  708.18 639.96 712.04 641.0 ;
      RECT  713.62 639.96 718.84 641.0 ;
      RECT  720.42 639.96 724.96 641.0 ;
      RECT  726.54 639.96 730.4 641.0 ;
      RECT  731.98 639.96 736.52 641.0 ;
      RECT  738.1 639.96 743.32 641.0 ;
      RECT  744.9 639.96 750.12 641.0 ;
      RECT  751.7 639.96 755.56 641.0 ;
      RECT  757.14 639.96 761.68 641.0 ;
      RECT  763.26 639.96 768.48 641.0 ;
      RECT  770.06 639.96 774.6 641.0 ;
      RECT  776.18 639.96 780.04 641.0 ;
      RECT  781.62 639.96 786.84 641.0 ;
      RECT  788.42 639.96 792.96 641.0 ;
      RECT  794.54 639.96 799.76 641.0 ;
      RECT  801.34 639.96 805.2 641.0 ;
      RECT  806.78 639.96 812.0 641.0 ;
      RECT  813.58 639.96 818.8 641.0 ;
      RECT  820.38 639.96 824.92 641.0 ;
      RECT  826.5 639.96 830.36 641.0 ;
      RECT  831.94 639.96 837.16 641.0 ;
      RECT  838.74 639.96 842.6 641.0 ;
      RECT  844.18 639.96 848.72 641.0 ;
      RECT  850.3 639.96 855.52 641.0 ;
      RECT  857.1 639.96 862.32 641.0 ;
      RECT  863.9 639.96 867.76 641.0 ;
      RECT  869.34 639.96 873.88 641.0 ;
      RECT  875.46 639.96 880.0 641.0 ;
      RECT  881.58 639.96 886.8 641.0 ;
      RECT  888.38 639.96 893.6 641.0 ;
      RECT  895.18 639.96 899.72 641.0 ;
      RECT  901.3 639.96 905.16 641.0 ;
      RECT  906.74 639.96 911.28 641.0 ;
      RECT  912.86 639.96 918.08 641.0 ;
      RECT  919.66 639.96 924.2 641.0 ;
      RECT  925.78 639.96 931.0 641.0 ;
      RECT  932.58 639.96 936.44 641.0 ;
      RECT  938.02 639.96 942.56 641.0 ;
      RECT  944.14 639.96 949.36 641.0 ;
      RECT  950.94 639.96 954.8 641.0 ;
      RECT  956.38 639.96 961.6 641.0 ;
      RECT  963.18 639.96 968.4 641.0 ;
      RECT  969.98 639.96 973.84 641.0 ;
      RECT  975.42 639.96 979.96 641.0 ;
      RECT  981.54 639.96 986.76 641.0 ;
      RECT  988.34 639.96 993.56 641.0 ;
      RECT  995.14 639.96 999.0 641.0 ;
      RECT  1000.58 639.96 1005.12 641.0 ;
      RECT  1006.7 639.96 1011.92 641.0 ;
      RECT  1013.5 639.96 1018.04 641.0 ;
      RECT  1019.62 639.96 1087.4 641.0 ;
      RECT  1088.98 1.66 1245.16 2.8 ;
      RECT  1088.98 2.8 1245.16 638.82 ;
      RECT  1088.98 638.82 1245.16 639.96 ;
      RECT  1245.16 1.66 1248.1 2.8 ;
      RECT  1245.16 638.82 1248.1 639.96 ;
      RECT  2.8 1.66 5.74 2.8 ;
      RECT  2.8 638.82 5.74 641.0 ;
      RECT  5.74 1.66 160.56 2.8 ;
      RECT  5.74 2.8 160.56 638.82 ;
      RECT  5.74 638.82 160.56 641.0 ;
      RECT  1110.06 0.62 1248.56 1.66 ;
      RECT  1220.22 639.96 1248.56 641.0 ;
      RECT  1248.1 1.66 1248.56 2.8 ;
      RECT  1248.1 2.8 1248.56 638.82 ;
      RECT  1248.1 638.82 1248.56 639.96 ;
      RECT  2.34 0.62 30.0 1.66 ;
      RECT  2.34 1.66 2.8 2.8 ;
      RECT  2.34 2.8 2.8 638.82 ;
      RECT  2.34 638.82 2.8 641.0 ;
   END
END    sky130_sram_1r1w_128x512_128
END    LIBRARY
