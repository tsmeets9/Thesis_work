module pytorch_mapping #(
  parameter int IO_DATA_WIDTH = 8,
  parameter int ACCUMULATION_WIDTH = 32
  )
  (
   input logic clk, 
   input logic CE,
   input logic [31:0] output_channel,
   input logic signed [ACCUMULATION_WIDTH-1:0] data_32b [0:15],
   output logic [IO_DATA_WIDTH-1:0] data_8b [0:15]
  );
  
  real scales [0:63];
  real biases [0:63];
  real interm;
  real interm2;

  initial begin

    interm = 0;
    scales[0] = 0.002669966248636571;
    scales[1] = 0.001285026212572898;
    scales[2] = 0.003335646230988762;
    scales[3] = 0.0015603260399029899;
    scales[4] = 0.0012292311904531683;
    scales[5] = 0.0017299280584317264;
    scales[6] = 0.0011421750282105847;
    scales[7] = 0.002278255156556215;
    scales[8] = 0.0020969203557169853;
    scales[9] = 0.0013154647735514756;
    scales[10] = 0.000993483645047032;
    scales[11] = 0.0031521873259591385;
    scales[12] = 0.0017990856190021325;
    scales[13] = 0.0015252230644664992;
    scales[14] = 0.0007723708381433357;
    scales[15] = 0.0010090796690468617;
    scales[16] = 0.0016940890865494204;
    scales[17] = 0.0013158821978776253;
    scales[18] = 0.0012806464332975648;
    scales[19] = 0.0010386160296056931;
    scales[20] = 0.0013965955465789566;
    scales[21] = 0.002266647505824001;
    scales[22] = 0.0035498453876658723;
    scales[23] = 0.0014903510342377637;
    scales[24] = 0.002243652185326115;
    scales[25] = 0.0011434730725452058;
    scales[26] = 0.002226981143580766;
    scales[27] = 0.0017085925152106767;
    scales[28] = 0.0016462649807731662;
    scales[29] = 0.002424689733403592;
    scales[30] = 0.0008702538405118084;
    scales[31] = 0.001563563101594208;
    scales[32] = 0.015652009155815046;
    scales[33] = 0.0010751888224891292;
    scales[34] = 0.0008734473933093274;
    scales[35] = 0.0036471887057169003;
    scales[36] = 0.0015335249094554505;
    scales[37] = 0.0008740687873291389;
    scales[38] = 0.0014377533936981986;
    scales[39] = 0.0012288213366745222;
    scales[40] = 0.001708925271229688;
    scales[41] = 0.005345158437513137;
    scales[42] = 0.002079191525748022;
    scales[43] = 0.002434429808382663;
    scales[44] = 0.0013832838265161204;
    scales[45] = 0.001203230449614119;
    scales[46] = 0.002037128345568688;
    scales[47] = 0.002193627921813281;
    scales[48] = 0.0019013012370051685;
    scales[49] = 0.0011524071017596062;
    scales[50] = 0.0010730233848497215;
    scales[51] = 0.00000008910621429590114;
    scales[52] = 0.002132520028683946;
    scales[53] = 0.0018194371650832818;
    scales[54] = 0.0011455762924666238;
    scales[55] = 0.0036482395325175224;
    scales[56] = 0.0005480913234295328;
    scales[57] = 0.0012104917359013609;
    scales[58] = 0.0019173346124044626;
    scales[59] = 0.002265671514320541;
    scales[60] = 0.0009994421880391332;
    scales[61] = 0.0008854554998991489;
    scales[62] = 0.0009803907747195028;
    scales[63] = 0.0006783627813566049;

    biases[0] = 69.89821;
    biases[1] = 9.303958;
    biases[2] = -70.41613;
    biases[3] = 41.598366;
    biases[4] = 39.27396;
    biases[5] = -7.776763;
    biases[6] = 14.435659;
    biases[7] = 42.92179;
    biases[8] = 16.934587;
    biases[9] = 25.446201;
    biases[10] = -8.922979;
    biases[11] = -48.583664;
    biases[12] = -13.226237;
    biases[13] = 52.761147;
    biases[14] = 28.21018;
    biases[15] = 31.738054;
    biases[16] = -33.789948;
    biases[17] = 37.246517;
    biases[18] = -21.34961;
    biases[19] = 2.9054353;
    biases[20] = -7.6019616;
    biases[21] = 64.83112;
    biases[22] = 49.16053;
    biases[23] = 6.6774926;
    biases[24] = -5.291203;
    biases[25] = -5.083957;
    biases[26] = -7.210429;
    biases[27] = -6.1439023;
    biases[28] = -10.790666;
    biases[29] = 42.533463;
    biases[30] = -1.8706831;
    biases[31] = -7.688503;
    biases[32] = -279.21967;
    biases[33] = -10.875337;
    biases[34] = 52.981358;
    biases[35] = 55.234272;
    biases[36] = -8.142929;
    biases[37] = 3.4470775;
    biases[38] = -12.946423;
    biases[39] = -24.106344;
    biases[40] = -15.014891;
    biases[41] = -21.718218;
    biases[42] = 48.500286;
    biases[43] = -18.765251;
    biases[44] = -7.3500037;
    biases[45] = 9.503984;
    biases[46] = 9.590292;
    biases[47] = -17.14792;
    biases[48] = -14.917725;
    biases[49] = 63.557495;
    biases[50] = -28.016172;
    biases[51] = -10.343923;
    biases[52] = 1.8994561;
    biases[53] = 47.442898;
    biases[54] = -18.429998;
    biases[55] = -86.702354;
    biases[56] = 19.106041;
    biases[57] = -19.54659;
    biases[58] = 7.91591;
    biases[59] = 27.45152;
    biases[60] = -20.015202;
    biases[61] = 24.400108;
    biases[62] = -18.593449;
    biases[63] = 15.419594;
  end 

  always @(posedge clk) begin
    if (CE) begin 
      for (int i=0; i<16; i++) begin 
        interm = scales[output_channel]*data_32b[i]+biases[output_channel];
        interm2 = (interm<0)? 0 : interm;
        data_8b[i] = $rtoi(interm2+0.5);
      end
    end
  end
endmodule

